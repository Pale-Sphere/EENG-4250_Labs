magic
tech scmos
timestamp 1758084387
<< nwell >>
rect 18 15 46 47
<< pwell >>
rect 6 -10 48 13
<< ntransistor >>
rect 24 -1 26 7
rect 34 -1 36 7
<< ptransistor >>
rect 26 32 34 34
rect 26 26 34 28
<< ndiffusion >>
rect 20 3 24 7
rect 22 -1 24 3
rect 26 3 28 7
rect 32 3 34 7
rect 26 -1 34 3
rect 36 3 40 7
rect 36 -1 38 3
<< pdiffusion >>
rect 26 35 28 38
rect 32 35 34 38
rect 26 34 34 35
rect 26 28 34 32
rect 26 25 34 26
rect 26 22 31 25
<< ndcontact >>
rect 18 -1 22 3
rect 28 3 32 7
rect 38 -1 42 3
<< pdcontact >>
rect 28 35 32 39
rect 31 21 35 25
<< psubstratepcontact >>
rect 10 -5 14 -1
<< nsubstratencontact >>
rect 39 35 43 39
<< polysilicon >>
rect 23 32 26 34
rect 34 32 42 34
rect 21 26 26 28
rect 34 26 37 28
rect 17 10 19 24
rect 40 18 42 32
rect 27 16 42 18
rect 36 10 38 16
rect 17 8 26 10
rect 24 7 26 8
rect 34 8 38 10
rect 34 7 36 8
rect 24 -4 26 -1
rect 34 -4 36 -1
<< polycontact >>
rect 17 24 21 28
rect 23 16 27 20
<< metal1 >>
rect 17 39 44 42
rect 32 13 35 21
rect 29 10 42 13
rect 29 7 32 10
rect 18 -5 21 -1
rect 39 -5 42 -1
rect 10 -8 42 -5
<< labels >>
rlabel metal1 18 -8 42 -5 5 GND!
rlabel metal1 17 39 42 42 1 Vdd!
rlabel polycontact 17 24 21 28 7 A
rlabel polycontact 23 16 27 20 7 B
rlabel metal1 38 10 42 13 3 out
<< end >>
