magic
tech scmos
timestamp 1758164354
<< polysilicon >>
rect 115 2 123 4
rect 115 -1 117 2
<< polycontact >>
rect 113 -5 117 -1
<< metal1 >>
rect -7 103 -3 107
rect -7 91 -3 95
rect -6 35 -2 39
rect -6 25 -2 29
rect 79 9 84 13
rect 79 1 89 5
rect 144 0 146 3
rect 108 -5 113 -2
rect -6 -34 -2 -30
rect -6 -46 -2 -42
rect -6 -102 -2 -98
rect -6 -115 -2 -111
<< m2contact >>
rect -3 102 3 107
rect -3 90 3 95
rect -2 34 4 39
rect -2 24 4 29
rect 73 9 79 14
rect 73 0 79 5
rect 146 -1 152 4
rect -2 -35 4 -30
rect -2 -47 4 -42
rect -2 -103 4 -98
rect -2 -115 4 -110
<< metal2 >>
rect 93 36 96 69
rect 76 33 96 36
rect 76 14 79 33
rect 68 0 73 3
rect 68 -34 71 0
rect 152 -1 155 4
rect 68 -37 96 -34
rect 93 -71 96 -37
use or4  or4_0
timestamp 1758161944
transform 1 0 50 0 1 52
box -50 -52 45 73
use or4  or4_1
timestamp 1758161944
transform 1 0 50 0 1 -85
box -50 -52 45 73
use nor2  nor2_0
timestamp 1758084387
transform 1 0 66 0 1 -15
box 6 -10 48 47
use inv  inv_0
timestamp 1758159428
transform 1 0 133 0 1 10
box -12 -35 15 19
<< labels >>
rlabel metal2 152 -1 155 4 3 out8
rlabel metal1 -7 103 -3 107 7 A
rlabel metal1 -7 91 -3 95 7 B
rlabel metal1 -6 35 -2 39 7 C
rlabel metal1 -6 25 -2 29 7 D
rlabel metal1 -6 -34 -2 -30 7 E
rlabel metal1 -6 -46 -2 -42 7 F
rlabel metal1 -6 -102 -2 -98 7 G
rlabel metal1 -6 -115 -2 -111 7 H
<< end >>
