magic
tech scmos
timestamp 1758066422
<< nwell >>
rect -12 -7 15 18
<< pwell >>
rect -12 -32 15 -8
<< ntransistor >>
rect 1 -21 9 -19
<< ptransistor >>
rect 1 4 8 6
<< ndiffusion >>
rect 1 -18 3 -14
rect 7 -18 9 -14
rect 1 -19 9 -18
rect 1 -22 9 -21
rect 1 -26 3 -22
rect 7 -26 9 -22
<< pdiffusion >>
rect 1 8 3 12
rect 7 8 8 12
rect 1 6 8 8
rect 1 3 8 4
rect 1 -1 3 3
rect 7 -1 8 3
<< ndcontact >>
rect 3 -18 7 -14
rect 3 -26 7 -22
<< pdcontact >>
rect 3 8 7 12
rect 3 -1 7 3
<< psubstratepcontact >>
rect -7 -28 -3 -24
<< nsubstratencontact >>
rect -7 11 -3 15
<< polysilicon >>
rect -10 4 1 6
rect 8 4 11 6
rect -10 -6 -8 4
rect -12 -8 -8 -6
rect -10 -19 -8 -8
rect -10 -21 1 -19
rect 9 -21 12 -19
<< metal1 >>
rect -6 15 6 17
rect -3 14 6 15
rect 3 12 6 14
rect 3 -7 6 -1
rect 3 -10 11 -7
rect 3 -14 6 -10
rect 3 -28 6 -26
rect -6 -31 6 -28
<< labels >>
rlabel metal1 8 -10 11 -7 1 out
rlabel metal1 4 15 5 16 5 Vdd!
rlabel metal1 4 -30 5 -29 1 GND!
rlabel polysilicon -12 -8 -10 -6 3 in
<< end >>
