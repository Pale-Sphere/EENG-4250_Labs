magic
tech scmos
timestamp 1758138774
<< nwell >>
rect -20 -4 31 27
<< pwell >>
rect -20 -22 31 -4
<< ntransistor >>
rect 3 -16 5 -10
rect 14 -16 16 -10
<< ptransistor >>
rect 3 2 5 9
rect 14 2 16 9
<< ndiffusion >>
rect -1 -11 3 -10
rect 0 -16 3 -11
rect 5 -16 14 -10
rect 16 -11 20 -10
rect 16 -16 19 -11
<< pdiffusion >>
rect -1 7 3 9
rect 0 2 3 7
rect 5 8 14 9
rect 5 3 7 8
rect 12 3 14 8
rect 5 2 14 3
rect 16 2 20 9
<< ndcontact >>
rect -5 -16 0 -11
rect 19 -16 24 -11
<< pdcontact >>
rect -5 2 0 7
rect 7 3 12 8
rect 20 2 25 7
<< psubstratepcontact >>
rect -15 -15 -10 -10
<< nsubstratencontact >>
rect -15 8 -10 13
<< polysilicon >>
rect 3 9 5 11
rect 14 9 16 11
rect 3 -10 5 2
rect 14 -10 16 2
rect 3 -19 5 -16
rect 14 -19 16 -16
<< polycontact >>
rect 1 11 6 16
rect 14 11 19 16
<< metal1 >>
rect -10 23 25 26
rect -10 7 -7 23
rect 1 16 4 20
rect 14 16 17 20
rect -10 4 -5 7
rect 22 7 25 23
rect 8 -1 11 3
rect 8 -4 23 -1
rect 20 -11 23 -4
rect -10 -15 -5 -12
<< labels >>
rlabel metal1 2 17 3 18 5 a
rlabel metal1 -9 5 -8 6 3 Vdd!
rlabel metal1 -9 -14 -8 -13 3 GND!
rlabel metal1 20 -4 22 -2 1 out
rlabel metal1 15 17 16 18 5 b
<< end >>
