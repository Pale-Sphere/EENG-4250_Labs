magic
tech scmos
timestamp 1757793793
<< pwell >>
rect 20 11 38 27
<< nwell >>
rect 20 -11 38 5
<< polysilicon >>
rect 21 18 25 20
rect 33 18 35 20
rect 21 9 23 18
rect 18 7 23 9
rect 21 -2 23 7
rect 21 -4 25 -2
rect 33 -4 35 -2
<< ndiffusion >>
rect 25 21 27 23
rect 31 21 33 23
rect 25 20 33 21
rect 25 17 33 18
rect 25 15 27 17
rect 31 15 33 17
<< pdiffusion >>
rect 25 -1 27 1
rect 31 -1 33 1
rect 25 -2 33 -1
rect 25 -5 33 -4
rect 25 -7 27 -5
rect 31 -7 33 -5
<< metal1 >>
rect 21 28 38 31
rect 28 25 31 28
rect 28 10 31 13
rect 28 7 34 10
rect 28 3 31 7
rect 28 -12 31 -9
rect 21 -15 38 -12
<< ntransistor >>
rect 25 18 33 20
<< ptransistor >>
rect 25 -4 33 -2
<< polycontact >>
rect 14 6 18 10
<< ndcontact >>
rect 27 21 31 25
rect 27 13 31 17
<< pdcontact >>
rect 27 -1 31 3
rect 27 -9 31 -5
<< labels >>
rlabel metal1 32 7 34 10 7 out
rlabel metal1 21 28 38 31 1 Vdd!
rlabel metal1 21 -15 38 -12 5 GND!
rlabel polysilicon 19 7 21 9 7 in
<< end >>
