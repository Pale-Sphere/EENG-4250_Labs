magic
tech scmos
timestamp 1758234173
<< metal1 >>
rect -52 51 -36 54
rect -52 42 -30 45
rect -4 44 17 47
rect -4 39 -1 44
rect -14 36 -1 39
rect 34 15 40 18
rect -51 -17 -36 -14
rect -51 -26 -29 -23
rect 25 -29 28 -12
rect -16 -32 28 -29
use nand2  nand2_0
timestamp 1758232332
transform 1 0 -9 0 1 3
box 10 -15 47 44
use nor2  nor2_0
timestamp 1758084387
transform 1 0 -53 0 1 26
box 6 -10 48 47
use nor2  nor2_1
timestamp 1758084387
transform 1 0 -53 0 1 -42
box 6 -10 48 47
<< labels >>
rlabel metal1 -50 -25 -50 -25 3 d
rlabel metal1 -50 -16 -50 -16 3 c
rlabel metal1 -51 52 -51 52 3 a
rlabel metal1 -51 43 -51 43 3 b
rlabel metal1 39 16 39 16 7 out4
<< end >>
