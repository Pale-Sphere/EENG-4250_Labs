magic
tech scmos
timestamp 1758159428
<< nwell >>
rect -12 -8 15 19
<< pwell >>
rect -12 -35 15 -8
<< ntransistor >>
rect 1 -23 9 -21
<< ptransistor >>
rect 1 5 8 7
<< ndiffusion >>
rect 1 -19 3 -14
rect 8 -19 9 -14
rect 1 -21 9 -19
rect 1 -24 9 -23
rect 1 -29 3 -24
rect 8 -29 9 -24
<< pdiffusion >>
rect 1 8 3 12
rect 1 7 8 8
rect 1 4 8 5
rect 1 -1 3 4
<< ndcontact >>
rect 3 -19 8 -14
rect 3 -29 8 -24
<< pdcontact >>
rect 3 8 8 13
rect 3 -1 8 4
<< psubstratepcontact >>
rect -8 -31 -3 -26
<< nsubstratencontact >>
rect -8 11 -3 16
<< polysilicon >>
rect -10 5 1 7
rect 8 5 11 7
rect -10 -6 -8 5
rect -12 -8 -8 -6
rect -10 -21 -8 -8
rect -10 -23 1 -21
rect 9 -23 12 -21
<< metal1 >>
rect -8 16 6 17
rect -3 14 6 16
rect 3 13 6 14
rect 3 -7 6 -1
rect 3 -10 11 -7
rect 3 -14 6 -10
rect 3 -31 6 -29
rect -6 -34 6 -31
<< labels >>
rlabel metal1 8 -10 11 -7 1 out
rlabel metal1 4 15 5 16 5 Vdd!
rlabel metal1 4 -33 5 -32 1 GND!
rlabel polysilicon -12 -8 -10 -6 3 in
<< end >>
